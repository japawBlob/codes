library verilog;
use verilog.vl_types.all;
entity majakEA_vlg_vec_tst is
end majakEA_vlg_vec_tst;
