library verilog;
use verilog.vl_types.all;
entity VGAgenerator_vlg_vec_tst is
end VGAgenerator_vlg_vec_tst;
