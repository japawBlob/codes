library verilog;
use verilog.vl_types.all;
entity NovaBlob_vlg_vec_tst is
end NovaBlob_vlg_vec_tst;
