library verilog;
use verilog.vl_types.all;
entity majakEA_vlg_check_tst is
    port(
        M               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end majakEA_vlg_check_tst;
